library	ieee;
use ieee.std_logic_1164.all;


entity test is
	
	
end entity;

architecture sim of test is

begin
	
	

end architecture;	