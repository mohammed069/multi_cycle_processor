library	ieee;
use ieee.std_logic_1164.all;


entity test is
	--generic
	
	--port 
	port(
	  x:in std_logic :='0';
	  y:out std_ulogic :='0'
	);
	
end entity;

architecture sim of test is
--declaration of architecture
begin
	--concurent statement
	

end architecture;	